`timescale 1ps / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/04/2021 10:54:15 AM
// Design Name: 
// Module Name: sra_control_ID_EX_stage
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sra_control_ID_EX_stage(
input signal_sra,input clock,output reg out_sra_control_reg);

always@(posedge clock)
out_sra_control_reg=signal_sra;
endmodule
